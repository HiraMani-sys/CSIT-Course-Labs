
LIBRARY ieee;
	USE ieee.std_logic_1164.ALL;

ENTITY NORGATE_HIRA IS
	PORT (
	A : IN STD_LOGIC;
	B : IN STD_LOGIC;
	C : OUT STD_LOGIC
	);
END NORGATE_HIRA;

ARCHITECTURE BEHAVIOUR OF NORGATE_HIRA IS
BEGIN
C <= A NOR B;
END BEHAVIOUR;
