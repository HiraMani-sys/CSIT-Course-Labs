
LIBRARY ieee;
	USE ieee.std_logic_1164.ALL;

ENTITY ANDGATE_HIRA IS
	PORT (
	A : IN STD_LOGIC;
	B : IN STD_LOGIC;
	C : OUT STD_LOGIC
	);
END ANDGATE_HIRA;

ARCHITECTURE BEHAVIOUR OF ANDGATE_HIRA IS
BEGIN
C <= A AND B;
END BEHAVIOUR;