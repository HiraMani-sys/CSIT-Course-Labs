
LIBRARY ieee;
	USE ieee.std_logic_1164.ALL;

ENTITY XORGATE_HIRA IS
	PORT (
	A : IN STD_LOGIC;
	B : IN STD_LOGIC;
	C : OUT STD_LOGIC
	);
END XORGATE_HIRA;

ARCHITECTURE BEHAVIOUR OF XORGATE_HIRA IS
BEGIN
C <= A XOR B;
END BEHAVIOUR;