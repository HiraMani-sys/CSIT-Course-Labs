
LIBRARY ieee;
	USE ieee.std_logic_1164.ALL;

ENTITY XNORGATE_HIRA IS
	PORT (
	A : IN STD_LOGIC;
	B : IN STD_LOGIC;
	C : OUT STD_LOGIC
	);
END XNORGATE_HIRA;

ARCHITECTURE BEHAVIOUR OF XNORGATE_HIRA IS
BEGIN
C <= A XNOR B;
END BEHAVIOUR;
