
LIBRARY ieee;
	USE ieee.std_logic_1164.ALL;

ENTITY NANDGATE_HIRA IS
	PORT (
	A : IN STD_LOGIC;
	B : IN STD_LOGIC;
	C : OUT STD_LOGIC
	);
END NANDGATE_HIRA;

ARCHITECTURE BEHAVIOUR OF NANDGATE_HIRA IS
BEGIN
C <= A NAND B;
END BEHAVIOUR;
